`include "define.h"

module memory_arbiter

endmodule


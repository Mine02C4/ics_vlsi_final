`include "define.h"

module fetcher
  (
    input [31:0] instr,
    output  nextstate
  );
  `include "parameter.h"

endmodule

